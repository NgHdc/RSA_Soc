`timescale 1ns / 1ps

//======================================================================
// Module: mod (Modular Reduction / Remainder)
// Computes R = a mod n (Remainder) and Q = a / n (Quotient)
// Note: Uses a basic restoring division algorithm approach.
//======================================================================
module mod #(
    parameter WIDTH = 19 // Default width, overridden during instantiation
) (
    input wire [WIDTH-1:0] a, // Dividend
    input wire [WIDTH-1:0] n, // Divisor (Modulus)
    output wire [WIDTH-1:0] R, // Remainder (a mod n)
    output wire [WIDTH-1:0] Q  // Quotient (a / n) - Often unused for modulo op
);

    // Internal registers for calculation
    reg [WIDTH-1:0] A_reg; // Holds quotient bits as they are determined
    reg [WIDTH-1:0] N_reg; // Latched divisor/modulus
    reg [WIDTH:0]   p_reg; // Partial remainder (needs one extra bit for subtraction)

    integer i;

    // Combinational logic block to perform division/modulo
    // Use always_comb in SystemVerilog for clarity, or always @(*) in Verilog-2001
    always @(*) begin
        A_reg = a; // Initialize quotient register (will be overwritten)
        N_reg = n; // Latch modulus
        p_reg = {{(WIDTH+1){1'b0}}}; // Initialize partial remainder to 0

        // Perform restoring division steps
        for (i = 0; i < WIDTH; i = i + 1) begin
            // 1. Shift left: Append next bit of dividend 'a' (from A_reg) to partial remainder 'p_reg'
            p_reg = {p_reg[WIDTH-1:0], A_reg[WIDTH-1]};

            // 2. Shift dividend (A_reg) left (conceptually, though we overwrite bits later)
            //    We overwrite A_reg[0] later, so only need to shift upper bits if required elsewhere.
            //    Let's prepare A_reg for quotient bit insertion:
            if (WIDTH > 1) begin
                 A_reg[WIDTH-1:1] = A_reg[WIDTH-2:0]; // Make space for quotient bit at A_reg[0]
            end

            // 3. Subtract divisor 'n' (N_reg) from partial remainder 'p_reg'
            //    Extend N_reg to WIDTH+1 bits for subtraction
            p_reg = p_reg - {1'b0, N_reg};

            // 4. Check sign bit (MSB of p_reg)
            if (p_reg[WIDTH] == 1'b1) begin // If result is negative (p < N originally)
                // Restore: Add N back
                p_reg = p_reg + {1'b0, N_reg};
                // Set quotient bit to 0
                A_reg[0] = 1'b0;
            end else begin // If result is non-negative (p >= N originally)
                // Keep subtraction result
                // Set quotient bit to 1
                A_reg[0] = 1'b1;
            end
        end
        // After the loop, p_reg holds the remainder and A_reg holds the quotient
    end

    // Assign outputs
    assign R = p_reg[WIDTH-1:0]; // Remainder is the final value in p_reg (lower WIDTH bits)
    assign Q = A_reg;           // Quotient is built in A_reg
endmodule

//======================================================================
// Module: mod_exp (Modular Exponentiation)
// Computes result = (base ^ exponent) mod modulo
// Uses the right-to-left binary method (square-and-multiply)
//======================================================================
module mod_exp #(
    parameter WIDTH = 32 // Base width (e.g., 32-bit RSA numbers might use WIDTH=1024)
                         // Note: Internal operations handle 2*WIDTH bits
) (
    input wire clk,
    input wire reset, // Active high asynchronous or synchronous reset
    input wire [WIDTH*2-1:0] base,
    input wire [WIDTH*2-1:0] modulo,
    input wire [WIDTH*2-1:0] exponent,
    output wire finish, // Goes high when computation is complete
    output wire [WIDTH*2-1:0] result // Final result of exponentiation
);

    // State machine definition
    localparam IDLE   = 2'd0; // Optional: Idle state before starting
    localparam UPDATE = 2'd1; // Calculation state
    localparam HOLD   = 2'd2; // Finished state

    // Internal registers
    reg [WIDTH*2-1:0] base_reg;     // Holds current base^(2^i) mod modulo
    reg [WIDTH*2-1:0] modulo_reg;   // Latched modulus
    reg [WIDTH*2-1:0] exponent_reg; // Holds remaining exponent bits
    reg [WIDTH*2-1:0] result_reg;   // Accumulates the result
    reg [1:0]         state;        // Current state of the FSM

    // Wires for intermediate calculations
    // Multiplication results need up to 2 * (operand width) = 4*WIDTH bits
    wire [WIDTH*4-1:0] result_mult_base_full;
    wire [WIDTH*4-1:0] base_squared_full;
    wire [WIDTH*2-1:0] result_next_mod; // Result after multiplying by base and taking modulo
    wire [WIDTH*2-1:0] base_next_mod;   // Result after squaring base and taking modulo

    // Assign outputs
    assign finish = (state == HOLD);
    assign result = result_reg;

    // Perform the multiplications
    assign result_mult_base_full = result_reg * base_reg;
    assign base_squared_full     = base_reg * base_reg;

    // Instantiate the 'mod' module for modular reduction
    // Instance 1: Calculate (base_reg * base_reg) mod modulo_reg
    mod #(
        .WIDTH(WIDTH*2) // Operands are WIDTH*2 bits
    ) base_sq_mod_inst (
        .a(base_squared_full[WIDTH*2-1:0]), // Input is the lower 2*WIDTH bits of the full product
        .n(modulo_reg),                     // Modulus
        .R(base_next_mod),                  // Result of modulo operation
        .Q()                                // Quotient not needed
    );

    // Instance 2: Calculate (result_reg * base_reg) mod modulo_reg
    mod #(
        .WIDTH(WIDTH*2) // Operands are WIDTH*2 bits
    ) res_mult_base_mod_inst (
        .a(result_mult_base_full[WIDTH*2-1:0]), // Input is the lower 2*WIDTH bits of the full product
        .n(modulo_reg),                         // Modulus
        .R(result_next_mod),                    // Result of modulo operation
        .Q()                                    // Quotient not needed
    );

    // State machine and register updates
    always @(posedge clk or posedge reset) begin // Use posedge reset if it's synchronous
        if (reset) begin
            // Reset state and registers
            state        <= IDLE; // Or UPDATE if calculation starts immediately
            base_reg     <= base; // Load initial base
            modulo_reg   <= modulo; // Load modulus
            exponent_reg <= exponent; // Load exponent
            // Initial result for square-and-multiply is 1
            result_reg   <= {{(WIDTH*2-1){1'b0}}, 1'b1};
        end else begin
            // State transitions and actions
            case (state)
                IDLE: begin
                    // Optional: Wait for a start signal or transition immediately
                    if (exponent != 0) begin // Start if exponent is non-zero
                       base_reg     <= base; // Load initial base
                       modulo_reg   <= modulo; // Load modulus
                       exponent_reg <= exponent; // Load exponent
                       result_reg   <= {{(WIDTH*2-1){1'b0}}, 1'b1}; // Initialize result
                       state        <= UPDATE;
                    end else begin
                       // If exponent is 0, result is 1 (already set)
                       base_reg     <= base;
                       modulo_reg   <= modulo;
                       exponent_reg <= exponent;
                       result_reg   <= {{(WIDTH*2-1){1'b0}}, 1'b1};
                       state        <= HOLD; // Go directly to HOLD
                    end
                end

                UPDATE: begin
                    if (exponent_reg != 0) begin
                        // If the current exponent bit (LSB) is 1
                        if (exponent_reg[0]) begin
                            result_reg <= result_next_mod; // result = (result * base) mod modulo
                        end else begin
                            // result_reg remains unchanged for this step
                        end

                        // Square the base: base = (base * base) mod modulo
                        base_reg <= base_next_mod;

                        // Shift exponent right: exponent = exponent >> 1
                        exponent_reg <= exponent_reg >> 1;

                        // Stay in UPDATE state
                        state <= UPDATE;
                    end else begin
                        // Exponent is 0, calculation finished
                        state <= HOLD;
                    end
                end

                HOLD: begin
                    // Remain in HOLD state, computation is finished
                    state <= HOLD;
                end

                default: begin
                    // Go to a safe state in case of an unexpected state value
                    state <= IDLE;
                end
            endcase
        end
    end
endmodule


//======================================================================
// Module: inverter (Modular Multiplicative Inverse)
// Computes d = e^-1 mod totient, where totient = (p-1)*(q-1)
// Also finds the smallest odd integer e > 1 such that gcd(e, totient) = 1
// Uses the Extended Euclidean Algorithm.
//======================================================================
module inverter #(
    parameter WIDTH = 32 // Width of primes p, q
                         // Totient and intermediate values use 2*WIDTH bits
) (
    input wire clk,
    input wire reset, // Active high reset
    input wire [WIDTH-1:0] p, // Prime p
    input wire [WIDTH-1:0] q, // Prime q
    output wire finish,       // Goes high when e and d are found
    output wire [WIDTH*2-1:0] e, // Public exponent (output)
    output wire [WIDTH*2-1:0] d  // Private exponent (output)
);

    // State machine definition
    localparam FIND_E   = 3'd0; // State to find a suitable 'e'
    localparam UPDATING = 3'd1; // State for Euclidean algorithm steps
    localparam CHECK    = 3'd2; // State to check GCD and finalize 'd'
    localparam HOLDING  = 3'd3; // State when finished

    // Internal registers
    reg [WIDTH*2-1:0] totient_reg; // Holds (p-1)*(q-1)
    reg [WIDTH*2-1:0] e_candidate; // Current 'e' being tested
    reg [WIDTH*2-1:0] a_reg;       // 'a' value in Euclidean algorithm (gcd(a,b))
    reg [WIDTH*2-1:0] b_reg;       // 'b' value in Euclidean algorithm (remainder)
    // Registers for Bezout coefficients (d = x*e + y*totient)
    // Need signed registers because intermediate values can be negative
    reg signed [WIDTH*2:0] x_prev; // Coefficient for 'a' (becomes 'd') - extra bit for sign
    reg signed [WIDTH*2:0] x_curr; // Coefficient for 'b' - extra bit for sign
    reg [2:0] state;               // FSM state

    // Wires
    wire [WIDTH*2-1:0] totient = (p-1)*(q-1); // Calculate Euler's totient
    wire [WIDTH*2-1:0] quotient;      // q = a / b from 'mod' module
    wire [WIDTH*2-1:0] remainder;     // r = a % b from 'mod' module (b_next)

    // Extended Euclidean Algorithm update step (signed arithmetic)
    // x_next = x_prev - quotient * x_curr
    wire signed [WIDTH*2+1:0] quotient_ext = $signed({1'b0, quotient}); // Extend quotient for wider mult
    wire signed [WIDTH*2+1:0] x_mult_q = $signed(x_curr) * quotient_ext; // Wider intermediate product
    wire signed [WIDTH*2+1:0] x_next = $signed(x_prev) - x_mult_q;

    // Instantiate the 'mod' module to calculate remainder and quotient
    mod #(
        .WIDTH(WIDTH*2) // Operating on totient-sized numbers
    ) gcd_step (
        .a(a_reg),      // Dividend (current GCD candidate)
        .n(b_reg),      // Divisor (current remainder)
        .R(remainder),  // Output: a mod b
        .Q(quotient)    // Output: a / b
    );

    // Assign outputs
    assign finish = (state == HOLDING);
    assign e = e_candidate; // Final chosen 'e'

    // --- FIX for vlog-13069: Break down complex assignment for 'd' ---
    // Intermediate wire for the adjusted 'd' value when x_prev is negative
    // Note: Addition result can require WIDTH*2+1 bits if there's a carry-out
    wire signed [WIDTH*2:0] d_adjusted_signed = $signed(x_prev) + $signed({1'b0, totient_reg});

    // Assign final 'd', selecting based on sign of x_prev and taking lower bits
    assign d = (x_prev[WIDTH*2] == 1'b1) // Check sign bit of x_prev
               ? d_adjusted_signed[WIDTH*2-1:0]  // If negative, use adjusted value (lower bits)
               : x_prev[WIDTH*2-1:0];           // If positive, use x_prev directly (lower bits)
    // --- End of fix ---

    // State machine and register updates
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= FIND_E;
            // Initialize first candidate e=3 (must be > 1 and odd)
            e_candidate <= {{(WIDTH*2-1){1'b0}}, 3'd3};
            totient_reg <= totient; // Latch totient
            // Initialize Euclidean algorithm registers for first 'e'
            a_reg <= totient; // Start with gcd(totient, e)
            b_reg <= {{(WIDTH*2-1){1'b0}}, 3'd3};
            // Initial Bezout coefficients for t in r = s*a + t*b (where a=totient, b=e)
            // Init: (r_prev, r_curr)=(a,b); (s_prev, s_curr)=(1,0); (t_prev, t_curr)=(0,1)
            x_prev <= $signed(1'b0); // t_prev = 0
            x_curr <= $signed(1'b1); // t_curr = 1

        end else begin
            case (state)
                FIND_E: begin
                    // Calculate totient (should be stable after reset if p,q are inputs)
                    totient_reg <= totient;
                    // Initialize for the current e_candidate
                    a_reg <= totient_reg; // Start with gcd(totient, e_candidate)
                    b_reg <= e_candidate;
                    x_prev <= $signed(1'b0); // Reset Bezout t_prev
                    x_curr <= $signed(1'b1); // Reset Bezout t_curr
                    state <= UPDATING;       // Start Euclidean algorithm
                end

                UPDATING: begin
                    // Perform one step of the Extended Euclidean Algorithm
                    if (b_reg != 0) begin // If remainder is not yet zero
                        a_reg <= b_reg;         // a = old b
                        b_reg <= remainder;     // b = old a mod old b
                        x_prev <= x_curr;       // Update Bezout coefficients
                        x_curr <= x_next[WIDTH*2:0]; // Use calculated next coefficient (lower WIDTH*2+1 bits)
                        state <= UPDATING;    // Continue algorithm
                    end else begin
                        // Remainder (b_reg) is zero, GCD is in a_reg
                        state <= CHECK;
                    end
                end

                CHECK: begin
                    // Check if GCD(totient, e) == 1 (stored in a_reg)
                    if (a_reg == 1) begin
                        // GCD is 1, found a valid 'e'. 'd' is calculated from x_prev.
                        state <= HOLDING;
                    end else begin
                        // GCD is not 1, this 'e' is not suitable. Try next odd 'e'.
                        e_candidate <= e_candidate + 2; // Increment e by 2
                        state <= FIND_E; // Restart the process for the new 'e'
                    end
                end

                HOLDING: begin
                    // Stay in HOLDING state, valid e and d found.
                    state <= HOLDING;
                end

                default: begin
                    state <= FIND_E; // Go to a safe state
                end
            endcase
        end
    end
endmodule


//======================================================================
// Module: control (Top-level RSA control logic)
// Coordinates key generation (inverter) and encryption/decryption (mod_exp)
//======================================================================
module control #(
    parameter WIDTH = 32 // Width for p, q, and base message size
                         // Internal operations use up to 2*WIDTH
) (
    input wire clk,
    input wire reset,         // Reset for inverter (key generation)
    input wire reset1,        // Reset for mod_exp (encrypt/decrypt operation)
    input wire [WIDTH-1:0] p, // Prime p input
    input wire [WIDTH-1:0] q, // Prime q input
    input wire encrypt_decrypt, // Control: 1 for encrypt (use e), 0 for decrypt (use d)
    input wire [WIDTH-1:0] msg_in, // Input message (plaintext/ciphertext)
    output wire [WIDTH*2-1:0] msg_out, // Output ciphertext/plaintext
    output wire mod_exp_finish       // Indicates completion of mod_exp
);

    // Wires connecting sub-modules
    wire inverter_finish;     // Signal from inverter when key parts (e, d) are ready
    wire [WIDTH*2-1:0] e;     // Public exponent from inverter
    wire [WIDTH*2-1:0] d;     // Private exponent from inverter
    wire [WIDTH*2-1:0] modulo; // n = p * q

    // Calculate modulo n = p * q
    assign modulo = p * q; // Direct multiplication

    // Select the exponent based on the mode (encrypt/decrypt)
    wire [WIDTH*2-1:0] exponent_selected;
    assign exponent_selected = encrypt_decrypt ? e : d;

    // Registers to stabilize inputs to mod_exp module
    reg [WIDTH*2-1:0] exp_reg; // Registered selected exponent
    reg [WIDTH*2-1:0] msg_reg; // Registered and zero-extended message
    reg [WIDTH*2-1:0] mod_reg; // Registered modulus

    // Register inputs for mod_exp on clock edge
    // Consider enabling updates based on inverter_finish or other control signals
    always @(posedge clk) begin
        // Example: Reset registers if either reset is active
        // Adjust reset condition as needed for your application
        if (reset || reset1) begin // Using OR condition for simplicity, adjust if needed
             exp_reg <= 0;
             msg_reg <= 0;
             mod_reg <= 0;
        end else begin
            // Latch values - perhaps only latch when inverter is finished?
            // Example: Latch continuously unless reset
            // if (inverter_finish) begin // Uncomment if latching should wait
                 exp_reg <= exponent_selected; // Latch the chosen exponent
                 mod_reg <= modulo;            // Latch the calculated modulus
                 // Latch and zero-extend the message input to match mod_exp base width
                 msg_reg <= {{(WIDTH){1'b0}}, msg_in};
            // end // Uncomment if latching should wait
        end
    end

    // Instantiate the inverter module to find e and d
    inverter #(
        .WIDTH(WIDTH) // Pass parameter value
    ) key_gen_inverter (
        .clk(clk),
        .reset(reset), // Use 'reset' for key generation
        .p(p),
        .q(q),
        .finish(inverter_finish), // Output: indicates e, d are ready
        .e(e),                 // Output: public exponent
        .d(d)                  // Output: private exponent
    );

    // Instantiate the modular exponentiation module for encryption/decryption
    mod_exp #(
        .WIDTH(WIDTH) // Pass parameter value
    ) encrypt_decrypt_mod_exp (
        .clk(clk),
        .reset(reset1),      // Use 'reset1' to start/reset encryption/decryption
        .base(msg_reg),       // Input: registered message (base for exponentiation)
        .modulo(mod_reg),    // Input: registered modulus n
        .exponent(exp_reg),  // Input: registered exponent (e or d)
        .finish(mod_exp_finish), // Output: indicates encryption/decryption is done
        .result(msg_out)      // Output: ciphertext or plaintext result
    );

endmodule
